--Memória ROM com 16 endereços de 18 bits
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity ROM is
    port(   clk: in std_logic;
            endereco : in unsigned(6 downto 0);
            dado: out unsigned(17 downto 0)
    );
end entity;
architecture a_ROM of ROM is
    type mem is array (0 to 127) of unsigned(17 downto 0);
    constant conteudo_rom : mem := (
        -- caso endereco => conteudo
        0 =>  "000000000000000000",
        1 =>  "000000000000000000",
        2 =>  "100000000000100000", -- LDA #32
        3 =>  "010100000000000010", -- STA 2
        4 =>  "100000000000000001", -- LDA 1 
        5 =>  "010100000000000001", -- STA 1
        6 =>  "011100000000000001", -- STOREMEM* reg1
        7 =>  "100100000000000001", -- ADD #1 + AC
        8 =>  "010000000000000010", -- CMP 2 ****
        9 =>  "110000001111110000", -- BRANCH -4
        10 => "000000000000000000", 
		11 => "100000000000000010", -- LDA #2
        12 => "010100000000000001", -- STA 1
        13 => "000100000000000001", -- ADD reg1
        14 => "101100000000000000", -- STOREMEM* 0
		15 => "010000000000100000", -- CMP 32
        16 => "110000001111101000", -- BRANCH -3
		17 => "000000000000000000", 
        18 => "100000000000000011", -- LDA #3               
        19 => "010100000000000001", -- STA 1            
        20 => "000100000000000001", -- ADD reg1                 
		21 => "101100000000000000", -- STOREMEM* 0              
        22 => "010000000000100000", -- CMP 32           
		23 => "110000001111101000", -- BRANCH -3            
        24 => "000000000000000000",
		25 => "100000000000000101", -- LDA #5
        26 => "010100000000000001", -- STA 1
		27 => "000100000000000001", -- ADD reg1
        28 => "101100000000000000", -- STOREMEM* 0
		29 => "010000000000100000", -- CMP 32 
        30 => "110000001111101000", -- BRANCH -3
		31 => "000000000000000000",
        32 => "100000000000000111", -- LDA #7
		33 => "010100000000000001", -- STA 1
        34 => "000100000000000001", -- ADD reg1
		35 => "101100000000000000", -- STOREMEM* 0
        36 => "010000000000100000", -- CMP 32
		37 => "110000001111101000", -- BRANCH -3
        38 => "000000000000000000",
		39 => "100000000000000010", -- LDA #2
        40 => "011100000000000011", -- LOADMEM* 3
        41 => "100100000000000001", -- ADD #1
        42 => "010000000000000010", -- CMP 2 
        43 => "110000001111101000", -- BRANCH -3
        44 => "000000000000000000",
        45 => "000000000000000000",
        46 => "000000000000000000",
        -- abaixo: casos omissos => (zero em todos os bits)
        others => (others=>'0')
    );
    begin
    process(clk)
        begin
            if(rising_edge(clk)) then
                dado <= conteudo_rom(to_integer(endereco));
            end if;
    end process;
end architecture;